//author:
//time  :
